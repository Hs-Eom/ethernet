`timescale 1ns / 1ps
module sw_axis
  #(
    // number of prefix/postfix characters
    parameter			      PREFIX_CHARS = 31,
    parameter			      POSTFIX_CHARS = 0,
    // those values
    parameter [(8*PREFIX_CHARS)-1:0]  PREFIX_STRING = "SWITCHES CHANGED! NEW VALUE: 0x",
    parameter [(8*POSTFIX_CHARS)-1:0] POSTFIX_STRING = "",
    // GPIO input width
    parameter			      GPIO_WIDTH = 2,
    // output axi bus width
    parameter			      AXI_OUT_WIDTH = 8,
    // Flag indicating if an additional two CRLF bytes must be added on the end
    // This creates a newline
    parameter			      INCLUDE_CRLF = 1,

    // convert the input string to ascii
    parameter			      ASCII_DATA = 1




    )
   ( 
     input			clk,
     input			reset_n,

     // input gpio
     input [GPIO_WIDTH-1:0]	gpio_in,
   
     // output axi master
     output [AXI_OUT_WIDTH-1:0]	m_axis_data,
     output			m_axis_valid,
     output			m_axis_last,
     output [11:0]		m_axis_tuser,
     input			m_axis_ready
   
     );

   // debounce gpio in
   logic [GPIO_WIDTH-1:0]	gpio_in_debounced;
   logic [GPIO_WIDTH-1:0]	gpio_in_debounced_z;


   debounce
     #(
       .DEBOUNCE_LENGTH(15),
       .NUM_PINS(GPIO_WIDTH)
       )
   debounce_i
     (
      .clk(clk),
      .reset_n(reset_n),
      .gpio_in(gpio_in),
      .gpio_out(gpio_in_debounced)
      );
   
   
   // Edge detect on gpio
   // This detects if *any* of the input pins (after debounce) changed
   logic			gpio_changed;
   
   always@(posedge clk)
     begin
        if (!reset_n) begin
           gpio_changed <= 0;
           gpio_in_debounced_z <= 0;
           
        end
        else begin
           gpio_in_debounced_z <= gpio_in_debounced;
           
           if (gpio_in_debounced != gpio_in_debounced_z) begin
              gpio_changed <= 1;
              
           end
           else begin
              gpio_changed <= 0;
              
           end
        end
     end


   typedef enum                     {IDLE, PREFIX, DATA, POSTFIX, WAIT}  state_type;
   state_type current_state = IDLE;
   state_type next_state    = IDLE;
   
   
   // If we enable INCLUDE_CRLF, the POSTFIX_CHARS and POSTFIX_STRING are extended by 2 bytes
   //기존 문자열에 \r\n을 추가하기 위해 2바이트 확장한거.
   localparam			    POSTFIX_CHARS_CR = POSTFIX_CHARS+2;
   localparam [(8*(POSTFIX_CHARS_CR))-1:0] POSTFIX_STRING_CR = {POSTFIX_STRING,16'h0A0D};
   localparam				   PREFIX_LENGTH = PREFIX_CHARS*8/AXI_OUT_WIDTH;
   localparam				   POSTFIX_LENGTH = INCLUDE_CRLF ? POSTFIX_CHARS_CR*8/AXI_OUT_WIDTH : POSTFIX_CHARS*8/AXI_OUT_WIDTH;

   localparam              ASCII_WIDTH = 4;
   localparam				   DATA_LENGTH = ASCII_WIDTH;//ASCII로 나타내면 4bytes필요함 ASCII말고 일반적인 데이터로 보낼려면 2bytes(16bit)면 충분

   localparam				   PACKET_PADDING = 5;//wait에서 잠시 쉬는시간
   

   logic [(8*PREFIX_LENGTH)-1:0]	   prefix_buffer;
   logic [(8*POSTFIX_LENGTH)-1:0]	   postfix_buffer;
   logic [(8*DATA_LENGTH)-1:0]		   data_buffer;
   
   logic				   fifo_full;

   // state dependant variables
   logic [AXI_OUT_WIDTH-1:0]		   axis_data;
   logic				   axis_valid;
   logic				   axis_ready;
   logic				   axis_last;
   logic [11:0]				   axis_user;
   // User contains total output length
   assign axis_user = PREFIX_LENGTH + DATA_LENGTH + POSTFIX_LENGTH;

   
		     
   // count the time spent in each state
   logic [31:0]				   state_counter;

   always @(posedge clk)
     begin
        if(!reset_n) begin
           state_counter  <= '0;

        end
        else begin
           if (current_state != next_state) begin
              state_counter  <= '0;

           end
           else begin
              // otherwise increment counter and shift buffer
              state_counter <= state_counter  + 'd1;
           end
        end
     end
   

   always @(*)
     begin
        next_state = current_state;
        case (current_state)
          IDLE   :
            begin
               if (gpio_changed & ~fifo_full & axis_ready) begin
                  if (PREFIX_LENGTH > 0) begin
                     next_state = PREFIX;
                  end
                  else begin
                     // No prefix, skip to data
                     next_state = DATA;
                     
                  end
               end 
            end
          PREFIX  :
            begin
               if (state_counter == PREFIX_LENGTH-1) begin
                  next_state = DATA;

               end
            end
          DATA  :
            begin
               if (state_counter == DATA_LENGTH-1) begin
                  if (POSTFIX_LENGTH > 0) begin
                     next_state = POSTFIX;

                  end
                  else begin
                     next_state = WAIT;

                  end
               end
            end
          POSTFIX  :
            begin
               if (state_counter == POSTFIX_LENGTH-1) begin
                  // no padding, 
                  next_state = WAIT;

               end
            end
          WAIT  :
            begin
               if (state_counter >= PACKET_PADDING-1) begin
                  next_state = IDLE;
                  
               end
            end
          default:
            next_state = current_state;
        endcase
     end
   
   
   always @(posedge clk)
     begin
        if(!reset_n) begin
           current_state <= IDLE;
        end
        else begin
           current_state <= next_state;
        end

     end

logic [31:0] gpio_ascii;
always@(*) begin   
   case(gpio_in_debounced_z)
      2'b00 : begin
         gpio_ascii[31 -: 8] = 8'h32; //2
         gpio_ascii[(31-8) -: 8] = 8'h62; //b
         gpio_ascii[(31-16) -: 8] = 8'd30; //0
         gpio_ascii[(31-24) -: 8] = 8'd30; //0
      end
      2'b01 : begin
         gpio_ascii[31 -: 8] = 8'h32; //2
         gpio_ascii[(31-8) -: 8] = 8'h62; //b
         gpio_ascii[(31-16) -: 8] = 8'd30; //0
         gpio_ascii[(31-24) -: 8] = 8'd31; //1
      end
      2'b10 : begin
         gpio_ascii[31 -: 8] = 8'h32; //2
         gpio_ascii[(31-8) -: 8] = 8'h62; //b
         gpio_ascii[(31-16) -: 8] = 8'd31; //1
         gpio_ascii[(31-24) -: 8] = 8'd30; //0
      end
      2'b11 : begin
         gpio_ascii[31 -: 8] = 8'h32; //2
         gpio_ascii[(31-8) -: 8] = 8'h62; //b
         gpio_ascii[(31-16) -: 8] = 8'd31; //1
         gpio_ascii[(31-24) -: 8] = 8'd31; //1
      end
      default : begin
         gpio_ascii[31 -: 8] = 8'h58; //X
         gpio_ascii[(31-8) -: 8] = 8'h58; //X
         gpio_ascii[(31-16) -: 8] = 8'd58; //X
         gpio_ascii[(31-24) -: 8] = 8'd58; //X
      end
   endcase
end

   // Load buffers
   always_ff@(posedge clk) begin
      if (!reset_n == 1) begin
         prefix_buffer <= 0;
         data_buffer   <= 0;
         postfix_buffer   <= 0;
         
      end
      else begin
         
         // prefix
         if (next_state == PREFIX && current_state != PREFIX) begin
            prefix_buffer   <= {<<8{PREFIX_STRING}};
            
         end
         // and data
         if (next_state == DATA && current_state != DATA) begin
            if (ASCII_DATA) begin
               data_buffer <= {<<8{gpio_ascii}}; 
            end
            else begin
               data_buffer <= {<<8{gpio_in_debounced_z}}; 
            end   
            
         end
         // and postfix
         if (next_state == POSTFIX && current_state != POSTFIX) begin
            postfix_buffer   <= {<<8{POSTFIX_STRING_CR}};
            
         end

         // shift out buffers
         if (current_state == PREFIX) begin
            prefix_buffer <= prefix_buffer >> AXI_OUT_WIDTH;
         end
         if (current_state == DATA) begin
            data_buffer <= data_buffer >> AXI_OUT_WIDTH;
         end
         if (current_state == POSTFIX) begin
            postfix_buffer <= postfix_buffer >> AXI_OUT_WIDTH;
         end
         
      end
   end

   // drive last on the cycle before we go into idle state
   assign axis_last = (next_state == WAIT & current_state != WAIT) ? 1 : 0;

   always @(*)
     begin
        case (current_state)
          IDLE   :
            begin
               axis_valid = 0;
               axis_data  = 0;
               
            end
          PREFIX  :
            begin
               axis_valid = 1;
               axis_data  = prefix_buffer[AXI_OUT_WIDTH-1:0];
               
            end
          DATA  :
            begin
               axis_valid = 1;
               axis_data  = data_buffer[AXI_OUT_WIDTH-1:0];
               
            end
          POSTFIX  :
            begin
               axis_valid = 1;
               axis_data  = postfix_buffer[AXI_OUT_WIDTH-1:0];
            end
          WAIT   :
            begin
               axis_valid = 0;
               axis_data  = 0;

            end
          default:
            begin
               axis_valid = 0;
               axis_data  = 0;

            end
        endcase
     end // always @ (*)
   
   
   axis_data_fifo_tuser axis_data_fifo_tuser 
     (
      .s_axis_aresetn(reset_n),          
      .s_axis_aclk(clk),                
      .s_axis_tvalid(axis_valid),        
      .s_axis_tready(axis_ready),        
      .s_axis_tdata(axis_data),          
      .s_axis_tlast(axis_last),          
      .s_axis_tuser(axis_user),          
      .m_axis_tvalid(m_axis_valid),      
      .m_axis_tready(m_axis_ready),      
      .m_axis_tdata(m_axis_data),        
      .m_axis_tlast(m_axis_last),        
      .m_axis_tuser(),               
      .axis_wr_data_count(),  
      .prog_full(fifo_full)              
      );

   assign m_axis_tuser = axis_user;

   
endmodule
